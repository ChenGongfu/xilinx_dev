`ifdef _COMMON_INCLUDE_VH_
`else
    `include "clogb2.v"
`endif 